module EPC(in, out);

	parameter n = 32;

	input  [n-1:0] in;
	output [n-1:0] out;

	assign out = in;

endmodule 